-- GENERATED WITH MATLAB...

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package GOLAY_SEQS_pkg is 

	 type type_a16x8std is array (0 to 16-1) of std_logic_vector(0 to 7);
 	 constant Ga128_1 : type_a16x8std := ( 
 	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "00110000",
	 	 	 	 "10101001",
	 	 	 	 "11000000",
	 	 	 	 "01011001",
	 	 	 	 "00110000",
	 	 	 	 "10101001",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "00110000",
	 	 	 	 "10101001",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "11001111",
	 	 	 	 "01010110"); 
 
	 constant Ga128_2 : type_a16x8std := ( 
 	 	 	 	 "01101010",
	 	 	 	 "11110011",
	 	 	 	 "01100101",
	 	 	 	 "11111100",
	 	 	 	 "10010101",
	 	 	 	 "00001100",
	 	 	 	 "01100101",
	 	 	 	 "11111100",
	 	 	 	 "01101010",
	 	 	 	 "11110011",
	 	 	 	 "01100101",
	 	 	 	 "11111100",
	 	 	 	 "01101010",
	 	 	 	 "11110011",
	 	 	 	 "10011010",
	 	 	 	 "00000011"); 
 
	 constant Ga128_3 : type_a16x8std := ( 
 	 	 	 	 "00110000",
	 	 	 	 "10101001",
	 	 	 	 "11000000",
	 	 	 	 "01011001",
	 	 	 	 "11001111",
	 	 	 	 "01010110",
	 	 	 	 "11000000",
	 	 	 	 "01011001",
	 	 	 	 "11001111",
	 	 	 	 "01010110",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "11001111",
	 	 	 	 "01010110",
	 	 	 	 "11000000",
	 	 	 	 "01011001"); 
 
	 constant Ga128_4 : type_a16x8std := ( 
 	 	 	 	 "01100101",
	 	 	 	 "11111100",
	 	 	 	 "10010101",
	 	 	 	 "00001100",
	 	 	 	 "10011010",
	 	 	 	 "00000011",
	 	 	 	 "10010101",
	 	 	 	 "00001100",
	 	 	 	 "10011010",
	 	 	 	 "00000011",
	 	 	 	 "01101010",
	 	 	 	 "11110011",
	 	 	 	 "10011010",
	 	 	 	 "00000011",
	 	 	 	 "10010101",
	 	 	 	 "00001100"); 
 
	 constant Gb128_1 : type_a16x8std := ( 
 	 	 	 	 "11000000",
	 	 	 	 "01011001",
	 	 	 	 "11001111",
	 	 	 	 "01010110",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "11001111",
	 	 	 	 "01010110",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "00110000",
	 	 	 	 "10101001",
	 	 	 	 "00111111",
	 	 	 	 "10100110",
	 	 	 	 "11001111",
	 	 	 	 "01010110"); 
 
	 constant Gb128_2 : type_a16x8std := ( 
 "10010101","00001100","10011010","00000011","01101010","11110011","10011010","00000011","01101010","11110011","01100101","11111100","01101010","11110011","10011010","00000011"); 
 
	 constant Gb128_3 : type_a16x8std := ( 
 "11001111","01010110","00111111","10100110","00110000","10101001","00111111","10100110","11001111","01010110","00111111","10100110","11001111","01010110","11000000","01011001"); 
 
	 constant Gb128_4 : type_a16x8std := ( 
 "10011010","00000011","01101010","11110011","01100101","11111100","01101010","11110011","10011010","00000011","01101010","11110011","10011010","00000011","10010101","00001100"); 
 
end GOLAY_SEQS_pkg; 
